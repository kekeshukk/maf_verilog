library verilog;
use verilog.vl_types.all;
entity First_one_2 is
    port(
        f_0             : in     vl_logic;
        f_1             : in     vl_logic;
        P               : out    vl_logic;
        V               : out    vl_logic
    );
end First_one_2;
