//暂时不要
module Transformer(
	input			[23:0]							iM_A,
	input			[23:0]							iM_B,
	input			[23:0]							iM_C,
	input			[13:0]							iE_A,
	input			[13:0]							iE_B,
	input			[13:0]							iE_C,
	output		[23:0]							M_A,
	output		[23:0]							M_B,
	output		[23:0]							M_C,
	output		[11:0]							M_A_H
);

endmodule