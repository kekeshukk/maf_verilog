library verilog;
use verilog.vl_types.all;
entity MAP_Top is
end MAP_Top;
